//  
// Copyright (c) 2023 Imperas Software Ltd., www.imperas.com  
//   
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0  
//  
// Licensed under the Apache License, Version 2.0 (the "License");  
// you may not use this file except in compliance with the License.  
// You may obtain a copy of the License at  
//  
//   http://www.apache.org/licenses/LICENSE-2.0  
//  
// Unless required by applicable law or agreed to in writing, software  
// distributed under the License is distributed on an "AS IS" BASIS,  
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,  
// either express or implied.  
//  
// See the License for the specific language governing permissions and  
// limitations under the License.  
//  
//  
 

typedef struct {
    string ins_str;
    ops_t ops[6];
    int hart;
    int issue;
    bit trap;
} ins_rv32i_t;


covergroup add_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add";
    
    cp_asm_count : coverpoint ins.ins_str == "add"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "GPR hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif

endgroup

covergroup addi_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add signed immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "addi"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup and_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "AND";
    
    cp_asm_count : coverpoint ins.ins_str == "and"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "GPR hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif

endgroup

covergroup andi_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "And signed immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "andi"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup auipc_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add upper immediate to PC";
    
    cp_asm_count : coverpoint ins.ins_str == "auipc"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup beq_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Equal";
    
    cp_asm_count : coverpoint ins.ins_str == "beq"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup bge_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Greater or Equal";
    
    cp_asm_count : coverpoint ins.ins_str == "bge"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup bgeu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Greater or Equal Unsigned";
    
    cp_asm_count : coverpoint ins.ins_str == "bgeu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup blt_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Less Than";
    
    cp_asm_count : coverpoint ins.ins_str == "blt"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup bltu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Less Than Unsigned";
    
    cp_asm_count : coverpoint ins.ins_str == "bltu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup bne_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Not Equal";
    
    cp_asm_count : coverpoint ins.ins_str == "bne"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_offset : coverpoint ins.ops[2].key.atohex() - get_pc(ins.hart, ins.issue, 0)  iff (ins.trap == 0 ) {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup jal_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Jump and Link";
    
    cp_asm_count : coverpoint ins.ins_str == "jal"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup jalr_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Jump and Link, register";
    
    cp_asm_count : coverpoint ins.ins_str == "jalr"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup lb_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Byte (8-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "lb"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory unaligned access";
    }
`endif

endgroup

covergroup lbu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Unsigned Byte (8-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "lbu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory unaligned access";
    }
`endif

endgroup

covergroup lh_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Half word (16-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "lh"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory unaligned access";
    }
`endif

endgroup

covergroup lhu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Unsigned Half word (16-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "lhu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory unaligned access";
    }
`endif

endgroup

covergroup lui_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Upper Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "lui"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup lw_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Word (32-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "lw"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "Memory unaligned access";
    }
`endif

endgroup

covergroup or_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "OR";
    
    cp_asm_count : coverpoint ins.ins_str == "or"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "GPR hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif

endgroup

covergroup ori_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Or signed immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "ori"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup sb_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Byte (8-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "sb"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup sh_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Half-word (16-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "sh"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup sll_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Left Logical";
    
    cp_asm_count : coverpoint ins.ins_str == "sll"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
`endif

endgroup

covergroup slli_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Left Logical Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "slli"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup slt_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less Than";
    
    cp_asm_count : coverpoint ins.ins_str == "slt"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
`endif

endgroup

covergroup slti_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less than Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "slti"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup sltiu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less than Immediate Unsigned";
    
    cp_asm_count : coverpoint ins.ins_str == "sltiu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup sltu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less Than Unsigned";
    
    cp_asm_count : coverpoint ins.ins_str == "sltu"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
`endif

endgroup

covergroup sra_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Arithmetic";
    
    cp_asm_count : coverpoint ins.ins_str == "sra"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
`endif

endgroup

covergroup srai_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Arithmetic Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "srai"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup srl_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Logical";
    
    cp_asm_count : coverpoint ins.ins_str == "srl"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
`endif

endgroup

covergroup srli_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Logical Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "srli"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup

covergroup sub_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Subtract";
    
    cp_asm_count : coverpoint ins.ins_str == "sub"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "GPR hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif

endgroup

covergroup sw_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Word (32-bit)";
    
    cp_asm_count : coverpoint ins.ins_str == "sw"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif

endgroup

covergroup xor_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Exlusive OR";
    
    cp_asm_count : coverpoint ins.ins_str == "xor"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) register assignment";
    }
    cp_rs2_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cmp_rs1_rs2_eq : coverpoint ins.ops[1].key == ins.ops[2].key  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rs1_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs2_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs2_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
    cr_rd_rs2 : cross cp_rd,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS2 register assignment";
    }
    cr_rd_rs1_rs2 : cross cp_rd,cp_rs1,cp_rs2  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD, RS1, and RS2 register assignment";
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 ) {
        option.comment = "GPR hazards";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif

endgroup

covergroup xori_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Exlusive-OR Immediate";
    
    cp_asm_count : coverpoint ins.ins_str == "xori"  iff (ins.trap == 0 ) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rd_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs1_sign : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint get_imm(ins.ops[2].key)  iff (ins.trap == 0 ) {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
    cp_rs1_maxvals : coverpoint unsigned'(get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER))  iff (ins.trap == 0 ) {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cmp_rd_rs1_eq : coverpoint ins.ops[0].key == ins.ops[1].key  iff (ins.trap == 0 ) {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.ops[0].key == "x0");
        bins x1  = {1} iff (ins.ops[0].key == "x1");
        bins x2  = {1} iff (ins.ops[0].key == "x2");
        bins x3  = {1} iff (ins.ops[0].key == "x3");
        bins x4  = {1} iff (ins.ops[0].key == "x4");
        bins x5  = {1} iff (ins.ops[0].key == "x5");
        bins x6  = {1} iff (ins.ops[0].key == "x6");
        bins x7  = {1} iff (ins.ops[0].key == "x7");
        bins x8  = {1} iff (ins.ops[0].key == "x8");
        bins x9  = {1} iff (ins.ops[0].key == "x9");
        bins x10  = {1} iff (ins.ops[0].key == "x10");
        bins x11  = {1} iff (ins.ops[0].key == "x11");
        bins x12  = {1} iff (ins.ops[0].key == "x12");
        bins x13  = {1} iff (ins.ops[0].key == "x13");
        bins x14  = {1} iff (ins.ops[0].key == "x14");
        bins x15  = {1} iff (ins.ops[0].key == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.ops[0].key == "x16");
        bins x17  = {1} iff (ins.ops[0].key == "x17");
        bins x18  = {1} iff (ins.ops[0].key == "x18");
        bins x19  = {1} iff (ins.ops[0].key == "x19");
        bins x20  = {1} iff (ins.ops[0].key == "x20");
        bins x21  = {1} iff (ins.ops[0].key == "x21");
        bins x22  = {1} iff (ins.ops[0].key == "x22");
        bins x23  = {1} iff (ins.ops[0].key == "x23");
        bins x24  = {1} iff (ins.ops[0].key == "x24");
        bins x25  = {1} iff (ins.ops[0].key == "x25");
        bins x26  = {1} iff (ins.ops[0].key == "x26");
        bins x27  = {1} iff (ins.ops[0].key == "x27");
        bins x28  = {1} iff (ins.ops[0].key == "x28");
        bins x29  = {1} iff (ins.ops[0].key == "x29");
        bins x30  = {1} iff (ins.ops[0].key == "x30");
        bins x31  = {1} iff (ins.ops[0].key == "x31");
`endif
    }
    cmp_rd_rs1_eqval : coverpoint get_gpr_val(ins.hart, ins.issue, ins.ops[0].key, `SAMPLE_AFTER) == get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, `SAMPLE_AFTER)  iff (ins.trap == 0 ) {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cr_rd_rs1 : cross cp_rd,cp_rs1  iff (ins.trap == 0 ) {
        option.comment = "Cross coverage of RD and RS1 register assignment";
    }
`endif

endgroup




function ins_rv32i_t get_rv32i_inst(bit trap, int hart, int issue, string disass); // break and move this first bit out
    string insbin, ins_str, op[6], key, val;
    ins_rv32i_t ins;
    int num, i, j;
    string s = disass;
    foreach (disass[c]) begin
        s[c] = (disass[c] == ",")? " " : disass[c];
    end
    ins.hart = hart;
    ins.issue = issue;
    ins.trap = trap;
    num = $sscanf (s, "%s %s %s %s %s %s %s %s", insbin, ins_str, op[0], op[1], op[2], op[3], op[4], op[5]);
    ins.ins_str = ins_str;
    for (i=0; i<num-2; i++) begin
        key = op[i];
        ins.ops[i].key=op[i]; // in case we dont update it as an indexed
        ins.ops[i].val=""; // not used
        for (j = 0; j < key.len(); j++) begin // if indexed addressing, convert offset(rs1) to op[i].key=rs1 op[i+1].key=offset
            if (key[j] == "(") begin
                ins.ops[i].key = key.substr(0,j-1); // offset
                ins.ops[i+1].key = key.substr(j+1,key.len()-2);
                i++; // step over +1
                //$display("indirect ins_str(%s) op[0](%0s).key(%s) op[1](%s).key(%s) op[2](%s).key(%s) op[3](%s).key(%s)", 
                //    ins_str, op[0], ins.ops[0].key, op[1], ins.ops[1].key, op[2], ins.ops[2].key, op[3], ins.ops[3].key);
                break;
            end
        end
    end
    for (i=0; i<num-2; i++) begin
        if (ins.ops[i].key[0] == "x") begin
            int idx = get_gpr_num(ins.ops[i].key);
            //$display("SAMPLE: %0s op[%0d]=%0s gpr(%0d)", ins_str,i, ins.ops[i].key, idx);
            if (idx < 0) begin
                ins.ops[i].val = ins.ops[i].key; // it is an immed already there
            end else begin
                ins.ops[i].val = string'(this.rvvi.x_wdata[hart][issue][idx]);
            end
        end else begin
            ins.ops[i].val = ins.ops[i].key;
        end       
    end
    return ins;
endfunction

function void rv32i_sample(string inst_name, bit trap, int hart, int issue, string disass);
    case (inst_name)
        "add"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        add_cg.sample(ins); 
                    end
        "addi"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        addi_cg.sample(ins); 
                    end
        "and"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        and_cg.sample(ins); 
                    end
        "andi"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        andi_cg.sample(ins); 
                    end
        "auipc"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        auipc_cg.sample(ins); 
                    end
        "beq"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        beq_cg.sample(ins); 
                    end
        "bge"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        bge_cg.sample(ins); 
                    end
        "bgeu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        bgeu_cg.sample(ins); 
                    end
        "blt"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        blt_cg.sample(ins); 
                    end
        "bltu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        bltu_cg.sample(ins); 
                    end
        "bne"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[1].key;
                        bne_cg.sample(ins); 
                    end
        "jal"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        jal_cg.sample(ins); 
                    end
        "jalr"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        jalr_cg.sample(ins); 
                    end
        "lb"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, 0) + get_imm(ins.ops[2].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_LOAD;
                        lb_cg.sample(ins); 
                    end
        "lbu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, 0) + get_imm(ins.ops[2].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_LOAD;
                        lbu_cg.sample(ins); 
                    end
        "lh"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, 0) + get_imm(ins.ops[2].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_LOAD;
                        lh_cg.sample(ins); 
                    end
        "lhu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, 0) + get_imm(ins.ops[2].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_LOAD;
                        lhu_cg.sample(ins); 
                    end
        "lui"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        lui_cg.sample(ins); 
                    end
        "lw"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[1].key, 0) + get_imm(ins.ops[2].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_LOAD;
                        lw_cg.sample(ins); 
                    end
        "or"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        or_cg.sample(ins); 
                    end
        "ori"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        ori_cg.sample(ins); 
                    end
        "sb"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[2].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, 0) + get_imm(ins.ops[1].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_STORE;
                        sb_cg.sample(ins); 
                    end
        "sh"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[2].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, 0) + get_imm(ins.ops[1].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_STORE;
                        sh_cg.sample(ins); 
                    end
        "sll"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        sll_cg.sample(ins); 
                    end
        "slli"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        slli_cg.sample(ins); 
                    end
        "slt"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        slt_cg.sample(ins); 
                    end
        "slti"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        slti_cg.sample(ins); 
                    end
        "sltiu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        sltiu_cg.sample(ins); 
                    end
        "sltu"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        sltu_cg.sample(ins); 
                    end
        "sra"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        sra_cg.sample(ins); 
                    end
        "srai"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        srai_cg.sample(ins); 
                    end
        "srl"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        srl_cg.sample(ins); 
                    end
        "srli"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        srli_cg.sample(ins); 
                    end
        "sub"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        sub_cg.sample(ins); 
                    end
        "sw"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[2].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].mem_addr = get_gpr_val(ins.hart, ins.issue, ins.ops[2].key, 0) + get_imm(ins.ops[1].val);
                        rvviDataQ[hart][issue][0].inst_category = INST_CAT_STORE;
                        sw_cg.sample(ins); 
                    end
        "xor"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        rvviDataQ[hart][issue][0].has_rs2 = 1;
                        rvviDataQ[hart][issue][0].rs2 = ins.ops[2].key;
                        xor_cg.sample(ins); 
                    end
        "xori"     : begin ins_rv32i_t ins = get_rv32i_inst(trap, hart, issue, disass); 
                        rvviDataQ[hart][issue][0].has_rd = 1;
                        rvviDataQ[hart][issue][0].rd = ins.ops[0].key;
                        rvviDataQ[hart][issue][0].has_rs1 = 1;
                        rvviDataQ[hart][issue][0].rs1 = ins.ops[1].key;
                        xori_cg.sample(ins); 
                    end
    endcase
endfunction


