//  
// Copyright (c) 2024 Imperas Software Ltd., www.imperas.com  
//   
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0  
//  
// Licensed under the Apache License, Version 2.0 (the "License");  
// you may not use this file except in compliance with the License.  
// You may obtain a copy of the License at  
//  
//   http://www.apache.org/licenses/LICENSE-2.0  
//  
// Unless required by applicable law or agreed to in writing, software  
// distributed under the License is distributed on an "AS IS" BASIS,  
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,  
// either express or implied.  
//  
// See the License for the specific language governing permissions and  
// limitations under the License.  
//  
//  
 


    add_cg = new(); add_cg.set_inst_name("obj_add");
    addi_cg = new(); addi_cg.set_inst_name("obj_addi");
    and_cg = new(); and_cg.set_inst_name("obj_and");
    andi_cg = new(); andi_cg.set_inst_name("obj_andi");
    auipc_cg = new(); auipc_cg.set_inst_name("obj_auipc");
    beq_cg = new(); beq_cg.set_inst_name("obj_beq");
    bge_cg = new(); bge_cg.set_inst_name("obj_bge");
    bgeu_cg = new(); bgeu_cg.set_inst_name("obj_bgeu");
    blt_cg = new(); blt_cg.set_inst_name("obj_blt");
    bltu_cg = new(); bltu_cg.set_inst_name("obj_bltu");
    bne_cg = new(); bne_cg.set_inst_name("obj_bne");
    jal_cg = new(); jal_cg.set_inst_name("obj_jal");
    jalr_cg = new(); jalr_cg.set_inst_name("obj_jalr");
    lb_cg = new(); lb_cg.set_inst_name("obj_lb");
    lbu_cg = new(); lbu_cg.set_inst_name("obj_lbu");
    lh_cg = new(); lh_cg.set_inst_name("obj_lh");
    lhu_cg = new(); lhu_cg.set_inst_name("obj_lhu");
    lui_cg = new(); lui_cg.set_inst_name("obj_lui");
    lw_cg = new(); lw_cg.set_inst_name("obj_lw");
    or_cg = new(); or_cg.set_inst_name("obj_or");
    ori_cg = new(); ori_cg.set_inst_name("obj_ori");
    sb_cg = new(); sb_cg.set_inst_name("obj_sb");
    sh_cg = new(); sh_cg.set_inst_name("obj_sh");
    sll_cg = new(); sll_cg.set_inst_name("obj_sll");
    slli_cg = new(); slli_cg.set_inst_name("obj_slli");
    slt_cg = new(); slt_cg.set_inst_name("obj_slt");
    slti_cg = new(); slti_cg.set_inst_name("obj_slti");
    sltiu_cg = new(); sltiu_cg.set_inst_name("obj_sltiu");
    sltu_cg = new(); sltu_cg.set_inst_name("obj_sltu");
    sra_cg = new(); sra_cg.set_inst_name("obj_sra");
    srai_cg = new(); srai_cg.set_inst_name("obj_srai");
    srl_cg = new(); srl_cg.set_inst_name("obj_srl");
    srli_cg = new(); srli_cg.set_inst_name("obj_srli");
    sub_cg = new(); sub_cg.set_inst_name("obj_sub");
    sw_cg = new(); sw_cg.set_inst_name("obj_sw");
    xor_cg = new(); xor_cg.set_inst_name("obj_xor");
    xori_cg = new(); xori_cg.set_inst_name("obj_xori");





