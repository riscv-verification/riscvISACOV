//
// Copyright (c) 2023 Imperas Software Ltd., www.imperas.com
// 
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    addi_cg = new(); addi_cg.set_inst_name("obj_addi");
    ori_cg = new(); ori_cg.set_inst_name("obj_ori");
    andi_cg = new(); andi_cg.set_inst_name("obj_andi");
    lui_cg = new(); lui_cg.set_inst_name("obj_lui");
    auipc_cg = new(); auipc_cg.set_inst_name("obj_auipc");
    jal_cg = new(); jal_cg.set_inst_name("obj_jal");
    jalr_cg = new(); jalr_cg.set_inst_name("obj_jalr");
    beq_cg = new(); beq_cg.set_inst_name("obj_beq");
    bne_cg = new(); bne_cg.set_inst_name("obj_bne");
    blt_cg = new(); blt_cg.set_inst_name("obj_blt");
    bge_cg = new(); bge_cg.set_inst_name("obj_bge");
    bltu_cg = new(); bltu_cg.set_inst_name("obj_bltu");
    bgeu_cg = new(); bgeu_cg.set_inst_name("obj_bgeu");
    lb_cg = new(); lb_cg.set_inst_name("obj_lb");
    lh_cg = new(); lh_cg.set_inst_name("obj_lh");
    lw_cg = new(); lw_cg.set_inst_name("obj_lw");
    lbu_cg = new(); lbu_cg.set_inst_name("obj_lbu");
    lhu_cg = new(); lhu_cg.set_inst_name("obj_lhu");
    sb_cg = new(); sb_cg.set_inst_name("obj_sb");
    sh_cg = new(); sh_cg.set_inst_name("obj_sh");
    sw_cg = new(); sw_cg.set_inst_name("obj_sw");
    slti_cg = new(); slti_cg.set_inst_name("obj_slti");
    sltiu_cg = new(); sltiu_cg.set_inst_name("obj_sltiu");
    xori_cg = new(); xori_cg.set_inst_name("obj_xori");
    slli_cg = new(); slli_cg.set_inst_name("obj_slli");
    srli_cg = new(); srli_cg.set_inst_name("obj_srli");
    srai_cg = new(); srai_cg.set_inst_name("obj_srai");
    add_cg = new(); add_cg.set_inst_name("obj_add");
    sub_cg = new(); sub_cg.set_inst_name("obj_sub");
    sll_cg = new(); sll_cg.set_inst_name("obj_sll");
    slt_cg = new(); slt_cg.set_inst_name("obj_slt");
    sltu_cg = new(); sltu_cg.set_inst_name("obj_sltu");
    xor_cg = new(); xor_cg.set_inst_name("obj_xor");
    srl_cg = new(); srl_cg.set_inst_name("obj_srl");
    sra_cg = new(); sra_cg.set_inst_name("obj_sra");
    or_cg = new(); or_cg.set_inst_name("obj_or");
    and_cg = new(); and_cg.set_inst_name("obj_and");


