//  
// Copyright (c) 2024 Imperas Software Ltd., www.imperas.com  
//   
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0  
//  
// Licensed under the Apache License, Version 2.0 (the "License");  
// you may not use this file except in compliance with the License.  
// You may obtain a copy of the License at  
//  
//   http://www.apache.org/licenses/LICENSE-2.0  
//  
// Unless required by applicable law or agreed to in writing, software  
// distributed under the License is distributed on an "AS IS" BASIS,  
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,  
// either express or implied.  
//  
// See the License for the specific language governing permissions and  
// limitations under the License.  
//  
//  
 



typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_rv32i_t;


covergroup add_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "add"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup addi_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add signed immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "addi"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup and_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "AND";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "and"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup andi_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "And signed immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "andi"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup auipc_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Add upper immediate to PC";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "auipc"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_zero : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        bins zero  = {0};
        bins nonzero  = default;
    }
`endif

endgroup

covergroup beq_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Equal";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "beq"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup bge_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Greater or Equal";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "bge"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup bgeu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Greater or Equal Unsigned";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "bgeu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup blt_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Less Than";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "blt"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup bltu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Less Than Unsigned";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "bltu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup bne_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Branch if Not Equal";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "bne"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_nord_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup jal_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Jump and Link";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "jal"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_zero : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        bins zero  = {0};
        bins nonzero  = default;
    }
`endif

endgroup

covergroup jalr_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Jump and Link, register";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "jalr"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup lb_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Byte (8-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lb"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup lbu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Unsigned Byte (8-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lbu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup lh_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Half word (16-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lh"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup lhu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Unsigned Half word (16-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lhu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup lui_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Upper Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lui"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_zero : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        bins zero  = {0};
        bins nonzero  = default;
    }
`endif

endgroup

covergroup lw_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Load Word (32-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "lw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup or_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "OR";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "or"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup ori_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Or signed immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "ori"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup sb_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Byte (8-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sb"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  {
        option.comment = "Memory unaligned access";
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup sh_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Half-word (16-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sh"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  {
        option.comment = "Memory unaligned access";
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup sll_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Left Logical";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sll"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup slli_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Left Logical Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "slli"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:31]};
    }
`endif

endgroup

covergroup slt_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less Than";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "slt"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_rd_boolean : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
`endif

endgroup

covergroup slti_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less than Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "slti"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_rd_boolean : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
`endif

endgroup

covergroup sltiu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less than Immediate Unsigned";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sltiu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_rd_boolean : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
`endif

endgroup

covergroup sltu_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Set if Less Than Unsigned";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sltu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_rd_boolean : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
`endif

endgroup

covergroup sra_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Arithmetic";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sra"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup srai_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Arithmetic Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "srai"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:31]};
    }
`endif

endgroup

covergroup srl_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Logical";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "srl"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup srli_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Shift Right Logical Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "srli"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif


`ifdef COVER_TYPE_VALUES
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:31]};
    }
`endif

endgroup

covergroup sub_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Subtract";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sub"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup sw_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Store Word (32-bit)";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "sw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_mem_unaligned : coverpoint is_unaligned_mem_access(ins.hart, ins.issue)  {
        option.comment = "Memory unaligned access";
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup xor_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Exlusive OR";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "xor"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
`endif


`ifdef COVER_TYPE_HAZARD
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs2_maxvals : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint ins.current.rd == ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2_eq : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2_eq : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup

covergroup xori_cg with function sample(ins_rv32i_t ins);
    option.per_instance = 1; 
    option.comment = "Exlusive-OR Immediate";
  

`ifdef COVER_TYPE_ASM_COUNT
    cp_asm_count : coverpoint ins.ins_str == "xori"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
`endif


`ifdef COVER_TYPE_ASSIGNMENTS
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) register assignment";
    }
`endif


`ifdef COVER_TYPE_EQUAL
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
`endif


`ifdef COVER_TYPE_MAXVALS
    cp_rd_maxvals : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
    cp_rs1_maxvals : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Max values";
        bins zeros  = {0};
        bins min  = {32'b10000000000000000000000000000000};
        bins max  = {32'b01111111111111111111111111111111};
        bins ones  = {32'b11111111111111111111111111111111};
        bins one  = {32'b00000000000000000000000000000001};
        bins minp1  = {32'b10000000000000000000000000000001};
    }
`endif


`ifdef COVER_TYPE_REG_COMPARE
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "Compare register assignment";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_eq : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
`endif


`ifdef COVER_TYPE_SIGNS
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins zero  = {0};
        bins pos  = {[1:$]};
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 (GPR) sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_imm : cross cp_rs1_sign,cp_imm_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm sign";
    }
`endif


`ifdef COVER_TYPE_TOGGLE
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0_1  = (32'b???????????????????????????????0 => 32'b???????????????????????????????1);
        wildcard bins bit_1_0_1  = (32'b??????????????????????????????0? => 32'b??????????????????????????????1?);
        wildcard bins bit_2_0_1  = (32'b?????????????????????????????0?? => 32'b?????????????????????????????1??);
        wildcard bins bit_3_0_1  = (32'b????????????????????????????0??? => 32'b????????????????????????????1???);
        wildcard bins bit_4_0_1  = (32'b???????????????????????????0???? => 32'b???????????????????????????1????);
        wildcard bins bit_5_0_1  = (32'b??????????????????????????0????? => 32'b??????????????????????????1?????);
        wildcard bins bit_6_0_1  = (32'b?????????????????????????0?????? => 32'b?????????????????????????1??????);
        wildcard bins bit_7_0_1  = (32'b????????????????????????0??????? => 32'b????????????????????????1???????);
        wildcard bins bit_8_0_1  = (32'b???????????????????????0???????? => 32'b???????????????????????1????????);
        wildcard bins bit_9_0_1  = (32'b??????????????????????0????????? => 32'b??????????????????????1?????????);
        wildcard bins bit_10_0_1  = (32'b?????????????????????0?????????? => 32'b?????????????????????1??????????);
        wildcard bins bit_11_0_1  = (32'b????????????????????0??????????? => 32'b????????????????????1???????????);
        wildcard bins bit_12_0_1  = (32'b???????????????????0???????????? => 32'b???????????????????1????????????);
        wildcard bins bit_13_0_1  = (32'b??????????????????0????????????? => 32'b??????????????????1?????????????);
        wildcard bins bit_14_0_1  = (32'b?????????????????0?????????????? => 32'b?????????????????1??????????????);
        wildcard bins bit_15_0_1  = (32'b????????????????0??????????????? => 32'b????????????????1???????????????);
        wildcard bins bit_16_0_1  = (32'b???????????????0???????????????? => 32'b???????????????1????????????????);
        wildcard bins bit_17_0_1  = (32'b??????????????0????????????????? => 32'b??????????????1?????????????????);
        wildcard bins bit_18_0_1  = (32'b?????????????0?????????????????? => 32'b?????????????1??????????????????);
        wildcard bins bit_19_0_1  = (32'b????????????0??????????????????? => 32'b????????????1???????????????????);
        wildcard bins bit_20_0_1  = (32'b???????????0???????????????????? => 32'b???????????1????????????????????);
        wildcard bins bit_21_0_1  = (32'b??????????0????????????????????? => 32'b??????????1?????????????????????);
        wildcard bins bit_22_0_1  = (32'b?????????0?????????????????????? => 32'b?????????1??????????????????????);
        wildcard bins bit_23_0_1  = (32'b????????0??????????????????????? => 32'b????????1???????????????????????);
        wildcard bins bit_24_0_1  = (32'b???????0???????????????????????? => 32'b???????1????????????????????????);
        wildcard bins bit_25_0_1  = (32'b??????0????????????????????????? => 32'b??????1?????????????????????????);
        wildcard bins bit_26_0_1  = (32'b?????0?????????????????????????? => 32'b?????1??????????????????????????);
        wildcard bins bit_27_0_1  = (32'b????0??????????????????????????? => 32'b????1???????????????????????????);
        wildcard bins bit_28_0_1  = (32'b???0???????????????????????????? => 32'b???1????????????????????????????);
        wildcard bins bit_29_0_1  = (32'b??0????????????????????????????? => 32'b??1?????????????????????????????);
        wildcard bins bit_30_0_1  = (32'b?0?????????????????????????????? => 32'b?1??????????????????????????????);
        wildcard bins bit_31_0_1  = (32'b0??????????????????????????????? => 32'b1???????????????????????????????);
        wildcard bins bit_0_1_0  = (32'b???????????????????????????????1 => 32'b???????????????????????????????0);
        wildcard bins bit_1_1_0  = (32'b??????????????????????????????1? => 32'b??????????????????????????????0?);
        wildcard bins bit_2_1_0  = (32'b?????????????????????????????1?? => 32'b?????????????????????????????0??);
        wildcard bins bit_3_1_0  = (32'b????????????????????????????1??? => 32'b????????????????????????????0???);
        wildcard bins bit_4_1_0  = (32'b???????????????????????????1???? => 32'b???????????????????????????0????);
        wildcard bins bit_5_1_0  = (32'b??????????????????????????1????? => 32'b??????????????????????????0?????);
        wildcard bins bit_6_1_0  = (32'b?????????????????????????1?????? => 32'b?????????????????????????0??????);
        wildcard bins bit_7_1_0  = (32'b????????????????????????1??????? => 32'b????????????????????????0???????);
        wildcard bins bit_8_1_0  = (32'b???????????????????????1???????? => 32'b???????????????????????0????????);
        wildcard bins bit_9_1_0  = (32'b??????????????????????1????????? => 32'b??????????????????????0?????????);
        wildcard bins bit_10_1_0  = (32'b?????????????????????1?????????? => 32'b?????????????????????0??????????);
        wildcard bins bit_11_1_0  = (32'b????????????????????1??????????? => 32'b????????????????????0???????????);
        wildcard bins bit_12_1_0  = (32'b???????????????????1???????????? => 32'b???????????????????0????????????);
        wildcard bins bit_13_1_0  = (32'b??????????????????1????????????? => 32'b??????????????????0?????????????);
        wildcard bins bit_14_1_0  = (32'b?????????????????1?????????????? => 32'b?????????????????0??????????????);
        wildcard bins bit_15_1_0  = (32'b????????????????1??????????????? => 32'b????????????????0???????????????);
        wildcard bins bit_16_1_0  = (32'b???????????????1???????????????? => 32'b???????????????0????????????????);
        wildcard bins bit_17_1_0  = (32'b??????????????1????????????????? => 32'b??????????????0?????????????????);
        wildcard bins bit_18_1_0  = (32'b?????????????1?????????????????? => 32'b?????????????0??????????????????);
        wildcard bins bit_19_1_0  = (32'b????????????1??????????????????? => 32'b????????????0???????????????????);
        wildcard bins bit_20_1_0  = (32'b???????????1???????????????????? => 32'b???????????0????????????????????);
        wildcard bins bit_21_1_0  = (32'b??????????1????????????????????? => 32'b??????????0?????????????????????);
        wildcard bins bit_22_1_0  = (32'b?????????1?????????????????????? => 32'b?????????0??????????????????????);
        wildcard bins bit_23_1_0  = (32'b????????1??????????????????????? => 32'b????????0???????????????????????);
        wildcard bins bit_24_1_0  = (32'b???????1???????????????????????? => 32'b???????0????????????????????????);
        wildcard bins bit_25_1_0  = (32'b??????1????????????????????????? => 32'b??????0?????????????????????????);
        wildcard bins bit_26_1_0  = (32'b?????1?????????????????????????? => 32'b?????0??????????????????????????);
        wildcard bins bit_27_1_0  = (32'b????1??????????????????????????? => 32'b????0???????????????????????????);
        wildcard bins bit_28_1_0  = (32'b???1???????????????????????????? => 32'b???0????????????????????????????);
        wildcard bins bit_29_1_0  = (32'b??1????????????????????????????? => 32'b??0?????????????????????????????);
        wildcard bins bit_30_1_0  = (32'b?1?????????????????????????????? => 32'b?0??????????????????????????????);
        wildcard bins bit_31_1_0  = (32'b1??????????????????????????????? => 32'b0???????????????????????????????);
    }
`endif

endgroup








function void rv32i_sample(int hart, int issue);
    ins_rv32i_t ins;

    case (traceDataQ[hart][issue][0].inst_name)
        "add"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            add_cg.sample(ins); 
        end
        "addi"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            addi_cg.sample(ins); 
        end
        "and"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            and_cg.sample(ins); 
        end
        "andi"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            andi_cg.sample(ins); 
        end
        "auipc"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            auipc_cg.sample(ins); 
        end
        "beq"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            beq_cg.sample(ins); 
        end
        "bge"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bge_cg.sample(ins); 
        end
        "bgeu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bgeu_cg.sample(ins); 
        end
        "blt"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            blt_cg.sample(ins); 
        end
        "bltu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bltu_cg.sample(ins); 
        end
        "bne"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bne_cg.sample(ins); 
        end
        "jal"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm_addr(1);
            jal_cg.sample(ins); 
        end
        "jalr"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm_addr(2);
            jalr_cg.sample(ins); 
        end
        "lb"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lb_cg.sample(ins); 
        end
        "lbu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lbu_cg.sample(ins); 
        end
        "lh"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lh_cg.sample(ins); 
        end
        "lhu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lhu_cg.sample(ins); 
        end
        "lui"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            lui_cg.sample(ins); 
        end
        "lw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lw_cg.sample(ins); 
        end
        "or"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            or_cg.sample(ins); 
        end
        "ori"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            ori_cg.sample(ins); 
        end
        "sb"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sb_cg.sample(ins); 
        end
        "sh"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sh_cg.sample(ins); 
        end
        "sll"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sll_cg.sample(ins); 
        end
        "slli"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            slli_cg.sample(ins); 
        end
        "slt"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            slt_cg.sample(ins); 
        end
        "slti"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            slti_cg.sample(ins); 
        end
        "sltiu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            sltiu_cg.sample(ins); 
        end
        "sltu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sltu_cg.sample(ins); 
        end
        "sra"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sra_cg.sample(ins); 
        end
        "srai"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            srai_cg.sample(ins); 
        end
        "srl"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            srl_cg.sample(ins); 
        end
        "srli"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            srli_cg.sample(ins); 
        end
        "sub"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sub_cg.sample(ins); 
        end
        "sw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sw_cg.sample(ins); 
        end
        "xor"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            xor_cg.sample(ins); 
        end
        "xori"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            xori_cg.sample(ins); 
        end
    endcase
endfunction







