//  
// Copyright (c) 2023 Imperas Software Ltd., www.imperas.com  
//   
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0  
//  
// Licensed under the Apache License, Version 2.0 (the "License");  
// you may not use this file except in compliance with the License.  
// You may obtain a copy of the License at  
//  
//   http://www.apache.org/licenses/LICENSE-2.0  
//  
// Unless required by applicable law or agreed to in writing, software  
// distributed under the License is distributed on an "AS IS" BASIS,  
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,  
// either express or implied.  
//  
// See the License for the specific language governing permissions and  
// limitations under the License.  
//  
//  
 
package RISCV_coverage_pkg;

import idvPkg::*;
import rvviApiPkg::*;

import idvApiPkg::*;

//`include "coverage/RISCV_coverage_global.svh"
`include "coverage/RISCV_coverage_common.svh"
`include "coverage/RISCV_trace_data.svh"

`include "coverage/RISCV_config_checks.svh"
`include "coverage/RISCV_instruction_base.svh"

`include "coverage/RISCV_coverage_base.svh"

endpackage

